
`include "Master.sv"
`include "Slave.sv"
`timescale 1ns/1ps

module test();

logic clk=0; // Clock which is sent from the testbench to the master.
logic reset; // Reset which is sent from the testbench to all the modules.
logic start; // This signals the master to start the transmission (also the master will read "masterDataToSend" in order to send it to the slave).
logic slaveSelect; // This tells the master which slave to transmit to. It should be read by the master when "start" becomes high.
logic [7:0] masterDataToSend; // What data should the master send to the slave during the transmission
logic [7:0] masterDataReceived; // What data did the master receive from the slave during the past transmission
logic [7:0] slaveDataToSend; // What data should the slave send to the master during the transmission
logic [7:0] slaveDataReceived; // What data did the slave receive from the master during the past transmission
logic SCLK; // The clock generated by the master for the transmission. The master uses the "clk" to generate this signal. Both the master and the slave can only use this signal for synchronizing the transmission. 
logic CS; // The chip select signal used by the master to select a slave. If a slave is selected, the master should set its corresponding CS to 0 (active low).

logic MOSI_0; // The data signals going from the master to the slave.
logic MOSI_1; 
logic MOSI_2; 
logic MOSI_3; 

logic MISO_0; // The data signals going from the slave to the master.
logic MISO_1;
logic MISO_2;
logic MISO_3;

// Here we create an instance of the master
Master m1(
	clk, reset,
	start, slaveSelect, masterDataToSend, masterDataReceived,
	SCLK, CS, MOSI_0, MOSI_1,  MOSI_2, MOSI_3, MISO_0, MISO_1, MISO_2, MISO_3);

// Here we create 1 instances of the slave which is flash
Slave flash(
	reset,
	slaveDataToSend, slaveDataReceived,
	SCLK, CS, MOSI_0, MOSI_1,  MOSI_2, MOSI_3, MISO_0, MISO_1, MISO_2, MISO_3);


always begin 
	#1 clk=~clk;
	   SCLK=clk;
end

initial begin
	
        reset = 0; // Set reset to 1 in order to reset all the modules
	start = 1;
	masterDataToSend = 8'hAB;
	slaveDataToSend = 8'hDE;
	slaveSelect=0;
	CS=0;
	#2 start=0;

	for (int i=0;i<16;i++) begin
		#1;
	end

	masterDataToSend = 8'h22;
	slaveDataToSend = 8'h33;
	start = 1;
	CS=0; //because my chip select was disabled
	#2 start=0;
	
	for (int i=0;i<16;i++) begin
		#1;
	end

$stop;
end

endmodule
